`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module encoder_4_2bitwise(
output [1:0]y,
input [3:0]I
   ); 
assign y[0]=I[1]|I[3];
assign y[1]=I[2]+I[3];
endmodule
