`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module Binary_Gray_conv_tb;
reg [3:0]B;
wire [3:0]G;
Binary_gray_conv u1(.G(G),.B(B));
initial
begin
B=4'b0111;#10;
B=4'b1110;#10;
B=4'b1000;#10;
B=4'b1011;#10;
$finish;
end
endmodule
