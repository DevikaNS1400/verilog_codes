`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module Encoder4_2_tb;
reg I0,I1,I2,I3;
wire A,B;
Encoder4_2 u1(.A(A),.B(B),.I0(I0),.I1(I1),.I2(I2),.I3(I3));
initial 
begin
I3=0;I2=0;I1=0;I0=0;#10;
I3=0;I2=0;I1=1;I0=0;#10;
I3=0;I2=1;I1=0;I0=0;#10;
I3=1;I2=0;I1=0;I0=0;#10;
$finish;
end
endmodule
