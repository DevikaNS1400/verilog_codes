`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module demux_2_1_bitwise_tb;
reg D,S;
wire A,B;
demux2_1bitwise u1(.A(A),.B(B),.D(D),.S(S));
 initial 
 begin
 D=1;S=0;#10;
 D=1;S=1;#10;
 D=0;S=1;#10;
 D=1;S=1;#10;
 $finish;
 end
endmodule
