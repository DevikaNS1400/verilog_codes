`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module gray2bin_tb;
reg [3:0]G;
wire [3:0]B;
gray2bin u1(.B(B),.G(G));
initial 
begin
G=4'b0011;#10;
G=4'b1010;#10;
G=4'b1001;#10;
G=4'b0110;#10;
G=4'b0111;#10;
G=4'b0101;#10;
G=4'b1011;#10;
G=4'b1110;#10;
$finish;
end
endmodule
