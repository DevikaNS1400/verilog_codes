`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module d_latch_tb();
reg D,en;
wire Q;
d_latch u1(.Q(Q),.D(D),.en(en));
initial begin
$monitor($time,"en=%d,D=%d,Q=%d",en,D,Q);
en=1'b0;D=1'b1;#10;
en=1'b1;D=1'b0;#10;
D=1'b1;#10;
D=1'b0;#10;
$finish;
end
endmodule
