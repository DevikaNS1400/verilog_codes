`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module mux2_1_tb;
reg A,B,S;
wire Y;
mux2_1bitwise u1(.Y(Y),.A(A),.B(B),.S(S));
initial 
begin
A=0;B=1;S=0;#10;
A=0;B=1;S=1;#10;
A=1;B=0;S=0;#10;
A=1;B=0;S=1;#10;
$finish;
end
endmodule
