`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module d_latch(
output reg Q,
input D,en
);
always@(en or D)begin
if(en==1)
Q<=D;
end
endmodule

