`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module comparator_1b(
output Y1,
output Y2,
output Y3,
input A,
input B
    );
 not g1(w1,A);
 not g2(w2,B);
 and g3(Y1,A,w2);//A>B
 xnor g4(Y2,A,B);//A=B
 and g5(Y3,w1,B);//A<B
endmodule
