`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module dff2tff_tb();
wire Q,Qn;
reg T,clk;
dff2tff u1(.Q(Q),.Qn(Qn),.T(T),.clk(clk));
always #5 clk=~clk;
initial begin
clk=1'b0;T=1'b0;#10;
T=1'b1;#15;
T=1'b0;#10;
T=1'b1;#10;
$finish;
end
endmodule
