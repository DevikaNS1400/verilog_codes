`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module even_parity_udm_tb;
reg A3,A2,A1,A0;
wire y;
even_parity_udm u1(.y(y),.A3(A3),.A2(A2),.A1(A1),.A0(A0));
initial
begin
A3=0;A2=0;A1=0;A0=0;#10;
A3=0;A2=0;A1=0;A0=1;#10;
A3=0;A2=0;A1=1;A0=0;#10;
A3=0;A2=0;A1=1;A0=1;#10;
A3=0;A2=1;A1=0;A0=0;#10;
A3=0;A2=1;A1=0;A0=1;#10;
A3=0;A2=1;A1=1;A0=0;#10;
A3=0;A2=1;A1=1;A0=1;#10;
A3=1;A2=0;A1=0;A0=0;#10;
A3=1;A2=0;A1=0;A0=1;#10;
A3=1;A2=0;A1=1;A0=0;#10;
A3=1;A2=0;A1=1;A0=1;#10;
A3=1;A2=1;A1=0;A0=0;#10;
A3=1;A2=1;A1=0;A0=1;#10;
A3=1;A2=1;A1=1;A0=0;#10;
A3=1;A2=1;A1=1;A0=1;#10;
$finish;
end
endmodule
