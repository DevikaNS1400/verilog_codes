`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module XOR_using_NAND(
output Y,
input A,
input B
    );
wire w1,w2,w3;
nand g1(w1,A,B);
nand g2(w2,A,w1);
nand g3(w3,B,w1);
nand g4(Y,w2,w3);
endmodule
