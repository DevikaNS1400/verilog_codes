`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module FA_Dataflow(
output S,
output c_out,
input A,
input B,
input C
   );
assign S=A^B^C;
assign c_out=(A&B)|C&(A^B);
endmodule
