`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module XOR_USING_NAND_tb;
reg A,B;
wire Y;
XOR_using_NAND u1(.Y(Y),.A(A),.B(B));
initial
begin
A=0;B=0;#10;
A=0;B=1;#10;
A=1;B=0;#10;
A=1;B=1;#10;
$finish;
end
endmodule
