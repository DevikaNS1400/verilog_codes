`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module decoder2to4 (
   output [3:0]I ,
    input[1:0]S
    );

    assign I[0] = ~S[1] & ~S[0];
    assign I[1] = ~S[1] &  S[0];
    assign I[2] =  S[1] & ~S[0];
    assign I[3] =  S[1] &  S[0];

endmodule

