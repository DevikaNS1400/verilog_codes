`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module D_flip_flop(
output reg Q,
input D,clk
    );
always@(posedge clk)
Q<=D;
endmodule
