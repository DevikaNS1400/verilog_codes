`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module sr_flipflop(
output reg Q,
output Qn,
input S,
input R,
input clk
    );
assign Qn=~Q;
always@(posedge clk)begin
case({S,R})
2'b00:Q<=Q;
2'b01:Q<=1'b0;
2'b10:Q<=1'b1;
2'b11:Q<=1'bx;
endcase 
end
endmodule
