`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module FUll_Sub_Dataflow(
output D,
output B_out,
input A,
input B,
input C
    );
    
assign D=A^B^C;
assign B_out=(~A&B)|(~A&C)|B&C;
endmodule
