`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module counter_tb();
wire [1:0]q;
reg clk;
counter1 u1(.q(q),.clk(clk));
always #5 clk=~clk;
initial begin
clk=0;#50;
$finish;
end
endmodule
