`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module comparator_1b_tb;
reg A,B;
wire Y1,Y2,Y3;
comparator_1b u1(.Y1(Y1),.Y2(Y2),.Y3(Y3),.A(A),.B(B));
initial
begin
A=0;B=0;#10;
A=0;B=1;#10;
A=1;B=0;#10;
A=1;B=1;#10;
$finish;
end
endmodule
