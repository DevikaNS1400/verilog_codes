`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module Encoder4_2(
output A,
output B,
input I0,
input I1,
input I2,
input I3);
assign A= I3|I2;
assign B=I1|I3;
endmodule
