`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module Decoder2_4_tb;
reg [1:0]S;
wire [3:0]I;
decoder2to4 u1(.S(S),.I(I));
initial
begin
S[1]=0;S[0]=0;#10;
S[1]=0;S[0]=1;#10;
S[1]=1;S[0]=0;#10;
S[1]=1;S[0]=1;#10;
$finish;
end
endmodule
