`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module sr_latch(
output Q,
output Q_bar,
input R,
input S
    );
nor g1(Q,Q_bar,R);
nor g2(Q_bar,Q,S);
endmodule
